magic
tech sky130A
timestamp 1642599340
<< mvnmos >>
rect -5 -10 45 90
rect 75 -10 125 90
rect 155 -10 205 90
rect 235 -10 285 90
rect 315 -10 365 90
rect 395 -10 445 90
rect 475 -10 525 90
rect 555 -10 605 90
<< mvndiff >>
rect -35 80 -5 90
rect -35 0 -29 80
rect -11 0 -5 80
rect -35 -10 -5 0
rect 45 80 75 90
rect 45 0 51 80
rect 69 0 75 80
rect 45 -10 75 0
rect 125 80 155 90
rect 125 0 131 80
rect 149 0 155 80
rect 125 -10 155 0
rect 205 80 235 90
rect 205 0 211 80
rect 229 0 235 80
rect 205 -10 235 0
rect 285 80 315 90
rect 285 0 291 80
rect 309 0 315 80
rect 285 -10 315 0
rect 365 80 395 90
rect 365 0 371 80
rect 389 0 395 80
rect 365 -10 395 0
rect 445 80 475 90
rect 445 0 451 80
rect 469 0 475 80
rect 445 -10 475 0
rect 525 80 555 90
rect 525 0 531 80
rect 549 0 555 80
rect 525 -10 555 0
rect 605 80 635 90
rect 605 0 611 80
rect 629 0 635 80
rect 605 -10 635 0
<< mvndiffc >>
rect -29 0 -11 80
rect 51 0 69 80
rect 131 0 149 80
rect 211 0 229 80
rect 291 0 309 80
rect 371 0 389 80
rect 451 0 469 80
rect 531 0 549 80
rect 611 0 629 80
<< mvpsubdiff >>
rect -120 160 -40 200
rect 640 160 720 200
rect -120 120 -80 160
rect 680 120 720 160
rect -120 -80 -80 -40
rect 680 -80 720 -40
rect -120 -120 -40 -80
rect 640 -120 720 -80
<< mvpsubdiffcont >>
rect -40 160 640 200
rect -120 -40 -80 120
rect 680 -40 720 120
rect -40 -120 640 -80
<< poly >>
rect -5 130 45 140
rect -5 110 10 130
rect 30 110 45 130
rect -5 90 45 110
rect 75 90 125 140
rect 155 90 205 140
rect 235 130 285 140
rect 235 110 250 130
rect 270 110 285 130
rect 235 90 285 110
rect 315 130 365 140
rect 315 110 330 130
rect 350 110 365 130
rect 315 90 365 110
rect 395 90 445 140
rect 475 90 525 140
rect 555 130 605 140
rect 555 110 570 130
rect 590 110 605 130
rect 555 90 605 110
rect -5 -60 45 -10
rect 75 -30 125 -10
rect 75 -50 90 -30
rect 110 -50 125 -30
rect 75 -60 125 -50
rect 155 -30 205 -10
rect 155 -50 170 -30
rect 190 -50 205 -30
rect 155 -60 205 -50
rect 235 -60 285 -10
rect 315 -60 365 -10
rect 395 -30 445 -10
rect 395 -50 410 -30
rect 430 -50 445 -30
rect 395 -60 445 -50
rect 475 -30 525 -10
rect 475 -50 490 -30
rect 510 -50 525 -30
rect 475 -60 525 -50
rect 555 -60 605 -10
<< polycont >>
rect 10 110 30 130
rect 250 110 270 130
rect 330 110 350 130
rect 570 110 590 130
rect 90 -50 110 -30
rect 170 -50 190 -30
rect 410 -50 430 -30
rect 490 -50 510 -30
<< locali >>
rect -120 190 -40 200
rect -120 170 -110 190
rect -90 170 -40 190
rect -120 160 -40 170
rect 640 190 720 200
rect 640 170 690 190
rect 710 170 720 190
rect 640 160 720 170
rect -120 120 -80 160
rect 0 110 10 130
rect 30 110 50 130
rect 70 110 80 130
rect 200 110 210 130
rect 230 110 250 130
rect 270 110 280 130
rect 320 110 330 130
rect 350 110 370 130
rect 390 110 400 130
rect 520 110 530 130
rect 550 110 570 130
rect 590 110 600 130
rect 680 120 720 160
rect -35 80 -5 90
rect -35 0 -30 80
rect -10 0 -5 80
rect -35 -10 -5 0
rect 45 80 75 90
rect 45 0 51 80
rect 69 0 75 80
rect 45 -10 75 0
rect 125 80 155 90
rect 125 0 130 80
rect 150 0 155 80
rect 125 -10 155 0
rect 205 80 235 90
rect 205 0 211 80
rect 229 0 235 80
rect 205 -10 235 0
rect 285 80 315 90
rect 285 0 290 80
rect 310 0 315 80
rect 285 -10 315 0
rect 365 80 395 90
rect 365 0 371 80
rect 389 0 395 80
rect 365 -10 395 0
rect 445 80 475 90
rect 445 0 450 80
rect 470 0 475 80
rect 445 -10 475 0
rect 525 80 555 90
rect 525 0 531 80
rect 549 0 555 80
rect 525 -10 555 0
rect 605 80 635 90
rect 605 0 610 80
rect 630 0 635 80
rect 605 -10 635 0
rect -120 -80 -80 -40
rect 70 -50 90 -30
rect 110 -50 120 -30
rect 160 -50 170 -30
rect 190 -50 210 -30
rect 390 -50 410 -30
rect 430 -50 440 -30
rect 480 -50 490 -30
rect 510 -50 530 -30
rect 680 -80 720 -40
rect -120 -90 -40 -80
rect -120 -110 -110 -90
rect -90 -110 -40 -90
rect -120 -120 -40 -110
rect 640 -90 720 -80
rect 640 -110 690 -90
rect 710 -110 720 -90
rect 640 -120 720 -110
<< viali >>
rect -110 170 -90 190
rect 690 170 710 190
rect 50 110 70 130
rect 210 110 230 130
rect 370 110 390 130
rect 530 110 550 130
rect -30 0 -29 80
rect -29 0 -11 80
rect -11 0 -10 80
rect 130 0 131 80
rect 131 0 149 80
rect 149 0 150 80
rect 290 0 291 80
rect 291 0 309 80
rect 309 0 310 80
rect 450 0 451 80
rect 451 0 469 80
rect 469 0 470 80
rect 610 0 611 80
rect 611 0 629 80
rect 629 0 630 80
rect 50 -50 70 -30
rect 210 -50 230 -30
rect 370 -50 390 -30
rect 530 -50 550 -30
rect -110 -110 -90 -90
rect 690 -110 710 -90
<< metal1 >>
rect -120 515 -80 520
rect -120 485 -115 515
rect -85 485 -80 515
rect -120 195 -80 485
rect 680 515 720 520
rect 680 485 685 515
rect 715 485 720 515
rect -120 165 -115 195
rect -85 165 -80 195
rect -120 -85 -80 165
rect -40 435 0 440
rect -40 405 -35 435
rect -5 405 0 435
rect -40 80 0 405
rect 280 435 320 440
rect 280 405 285 435
rect 315 405 320 435
rect 40 355 80 360
rect 40 325 45 355
rect 75 325 80 355
rect 40 130 80 325
rect 200 355 240 360
rect 200 325 205 355
rect 235 325 240 355
rect 40 110 50 130
rect 70 110 80 130
rect 40 100 80 110
rect 120 275 160 280
rect 120 245 125 275
rect 155 245 160 275
rect -40 0 -30 80
rect -10 0 0 80
rect -40 -10 0 0
rect 120 80 160 245
rect 200 130 240 325
rect 200 110 210 130
rect 230 110 240 130
rect 200 100 240 110
rect 120 0 130 80
rect 150 0 160 80
rect 120 -10 160 0
rect 280 80 320 405
rect 600 435 640 440
rect 600 405 605 435
rect 635 405 640 435
rect 360 355 400 360
rect 360 325 365 355
rect 395 325 400 355
rect 360 130 400 325
rect 520 355 560 360
rect 520 325 525 355
rect 555 325 560 355
rect 360 110 370 130
rect 390 110 400 130
rect 360 100 400 110
rect 440 275 480 280
rect 440 245 445 275
rect 475 245 480 275
rect 280 0 290 80
rect 310 0 320 80
rect 280 -10 320 0
rect 440 80 480 245
rect 520 130 560 325
rect 520 110 530 130
rect 550 110 560 130
rect 520 100 560 110
rect 440 0 450 80
rect 470 0 480 80
rect 440 -10 480 0
rect 600 80 640 405
rect 600 0 610 80
rect 630 0 640 80
rect 600 -10 640 0
rect 680 195 720 485
rect 680 165 685 195
rect 715 165 720 195
rect -120 -115 -115 -85
rect -85 -115 -80 -85
rect -120 -485 -80 -115
rect 40 -30 80 -20
rect 40 -50 50 -30
rect 70 -50 80 -30
rect 40 -165 80 -50
rect 40 -195 45 -165
rect 75 -195 80 -165
rect 40 -200 80 -195
rect 200 -30 240 -20
rect 200 -50 210 -30
rect 230 -50 240 -30
rect 200 -245 240 -50
rect 200 -275 205 -245
rect 235 -275 240 -245
rect 200 -280 240 -275
rect 360 -30 400 -20
rect 360 -50 370 -30
rect 390 -50 400 -30
rect 360 -325 400 -50
rect 360 -355 365 -325
rect 395 -355 400 -325
rect 360 -360 400 -355
rect 520 -30 560 -20
rect 520 -50 530 -30
rect 550 -50 560 -30
rect 520 -405 560 -50
rect 520 -435 525 -405
rect 555 -435 560 -405
rect 520 -440 560 -435
rect 680 -85 720 165
rect 680 -115 685 -85
rect 715 -115 720 -85
rect -120 -515 -115 -485
rect -85 -515 -80 -485
rect -120 -520 -80 -515
rect 680 -485 720 -115
rect 680 -515 685 -485
rect 715 -515 720 -485
rect 680 -520 720 -515
<< via1 >>
rect -115 485 -85 515
rect 685 485 715 515
rect -115 190 -85 195
rect -115 170 -110 190
rect -110 170 -90 190
rect -90 170 -85 190
rect -115 165 -85 170
rect -35 405 -5 435
rect 285 405 315 435
rect 45 325 75 355
rect 205 325 235 355
rect 125 245 155 275
rect 605 405 635 435
rect 365 325 395 355
rect 525 325 555 355
rect 445 245 475 275
rect 685 190 715 195
rect 685 170 690 190
rect 690 170 710 190
rect 710 170 715 190
rect 685 165 715 170
rect -115 -90 -85 -85
rect -115 -110 -110 -90
rect -110 -110 -90 -90
rect -90 -110 -85 -90
rect -115 -115 -85 -110
rect 45 -195 75 -165
rect 205 -275 235 -245
rect 365 -355 395 -325
rect 525 -435 555 -405
rect 685 -90 715 -85
rect 685 -110 690 -90
rect 690 -110 710 -90
rect 710 -110 715 -90
rect 685 -115 715 -110
rect -115 -515 -85 -485
rect 685 -515 715 -485
<< metal2 >>
rect -120 515 720 520
rect -120 485 -115 515
rect -85 485 685 515
rect 715 485 720 515
rect -120 480 720 485
rect -120 435 720 440
rect -120 405 -35 435
rect -5 405 285 435
rect 315 405 605 435
rect 635 405 720 435
rect -120 400 720 405
rect -120 355 720 360
rect -120 325 45 355
rect 75 325 205 355
rect 235 325 365 355
rect 395 325 525 355
rect 555 325 720 355
rect -120 320 720 325
rect -120 275 720 280
rect -120 245 125 275
rect 155 245 445 275
rect 475 245 720 275
rect -120 240 720 245
rect -120 195 720 200
rect -120 165 -115 195
rect -85 165 685 195
rect 715 165 720 195
rect -120 160 720 165
rect -120 -85 720 -80
rect -120 -115 -115 -85
rect -85 -115 685 -85
rect 715 -115 720 -85
rect -120 -120 720 -115
rect -120 -165 720 -160
rect -120 -195 45 -165
rect 75 -195 720 -165
rect -120 -200 720 -195
rect -120 -245 720 -240
rect -120 -275 205 -245
rect 235 -275 720 -245
rect -120 -280 720 -275
rect -120 -325 720 -320
rect -120 -355 365 -325
rect 395 -355 720 -325
rect -120 -360 720 -355
rect -120 -405 720 -400
rect -120 -435 525 -405
rect 555 -435 720 -405
rect -120 -440 720 -435
rect -120 -485 720 -480
rect -120 -515 -115 -485
rect -85 -515 685 -485
rect 715 -515 720 -485
rect -120 -520 720 -515
<< labels >>
rlabel metal2 -120 400 -80 440 0 D
port 1 nsew
rlabel metal2 -120 320 -80 360 0 G
port 2 nsew
rlabel metal2 -120 240 -80 280 0 S
port 3 nsew
rlabel metal2 -120 160 -80 200 0 VSS
port 4 nsew
rlabel metal2 680 -200 720 -160 0 A1
port 5 nsew
rlabel metal2 680 -280 720 -240 0 A2
port 6 nsew
rlabel metal2 680 -360 720 -320 0 A3
port 7 nsew
rlabel metal2 680 -440 720 -400 0 A4
port 8 nsew
rlabel locali 50 30 70 50 0 B1
rlabel locali 210 30 230 50 0 B2
rlabel locali 370 30 390 50 0 B3
rlabel locali 530 30 550 50 0 B4
<< end >>
