* NGSPICE file created from prognmos.ext - technology: sky130A

.subckt prognmos D G S VSS A1 A2 A3 A4
X0 S A1 B1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
X1 B3 G D VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=2.25e+11p ps=1.95e+06u w=1e+06u l=500000u
X2 B1 G D VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=2.25e+11p ps=1.95e+06u w=1e+06u l=500000u
X3 B2 A2 S VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
X4 D G B4 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.25e+11p pd=1.95e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
X5 S A3 B3 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
X6 D G B2 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.25e+11p pd=1.95e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
X7 B4 A4 S VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.5e+11p pd=1.3e+06u as=1.5e+11p ps=1.3e+06u w=1e+06u l=500000u
.ends

