magic
tech sky130A
timestamp 1642601396
<< metal2 >>
rect -400 4435 -360 4440
rect -400 4405 -395 4435
rect -365 4405 -360 4435
rect -400 4355 -360 4405
rect -400 4325 -395 4355
rect -365 4325 -360 4355
rect -400 4320 -360 4325
rect -320 4435 -280 4440
rect -320 4405 -315 4435
rect -285 4405 -280 4435
rect -320 4355 -280 4405
rect -320 4325 -315 4355
rect -285 4325 -280 4355
rect -320 4320 -280 4325
rect 880 4435 920 4440
rect 880 4405 885 4435
rect 915 4405 920 4435
rect 880 4355 920 4405
rect 880 4325 885 4355
rect 915 4325 920 4355
rect 880 4320 920 4325
rect 960 4435 1000 4440
rect 960 4405 965 4435
rect 995 4405 1000 4435
rect 960 4355 1000 4405
rect 960 4325 965 4355
rect 995 4325 1000 4355
rect 960 4320 1000 4325
rect 1040 4435 1080 4440
rect 1040 4405 1045 4435
rect 1075 4405 1080 4435
rect 1040 4355 1080 4405
rect 1040 4325 1045 4355
rect 1075 4325 1080 4355
rect 1040 4320 1080 4325
rect 1120 4435 1160 4440
rect 1120 4405 1125 4435
rect 1155 4405 1160 4435
rect 1120 4355 1160 4405
rect 1120 4325 1125 4355
rect 1155 4325 1160 4355
rect 1120 4320 1160 4325
rect 1200 4435 1240 4440
rect 1200 4405 1205 4435
rect 1235 4405 1240 4435
rect 1200 4355 1240 4405
rect 1200 4325 1205 4355
rect 1235 4325 1240 4355
rect 1200 4320 1240 4325
rect 1280 4435 1320 4440
rect 1280 4405 1285 4435
rect 1315 4405 1320 4435
rect 1280 4355 1320 4405
rect 1280 4325 1285 4355
rect 1315 4325 1320 4355
rect 1280 4320 1320 4325
rect 1360 4435 1400 4440
rect 1360 4405 1365 4435
rect 1395 4405 1400 4435
rect 1360 4355 1400 4405
rect 1360 4325 1365 4355
rect 1395 4325 1400 4355
rect 1360 4320 1400 4325
rect 1440 4435 1480 4440
rect 1440 4405 1445 4435
rect 1475 4405 1480 4435
rect 1440 4355 1480 4405
rect 1440 4325 1445 4355
rect 1475 4325 1480 4355
rect 1440 4320 1480 4325
rect -400 4275 0 4280
rect -400 4245 -75 4275
rect -45 4245 0 4275
rect -400 4240 0 4245
rect -400 4195 0 4200
rect -400 4165 -395 4195
rect -365 4165 0 4195
rect -400 4160 0 4165
rect -400 4115 0 4120
rect -400 4085 -395 4115
rect -365 4085 0 4115
rect -400 4080 0 4085
rect -240 4035 0 4040
rect -240 4005 -235 4035
rect -205 4005 0 4035
rect -240 4000 0 4005
rect -80 3955 0 3960
rect -80 3925 -75 3955
rect -45 3925 0 3955
rect -80 3920 0 3925
rect -80 3675 0 3680
rect -80 3645 -75 3675
rect -45 3645 0 3675
rect -80 3640 0 3645
rect 840 3595 920 3600
rect 840 3565 885 3595
rect 915 3565 920 3595
rect 840 3560 920 3565
rect 840 3515 1000 3520
rect 840 3485 965 3515
rect 995 3485 1000 3515
rect 840 3480 1000 3485
rect 840 3435 1080 3440
rect 840 3405 1045 3435
rect 1075 3405 1080 3435
rect 840 3400 1080 3405
rect 840 3355 1160 3360
rect 840 3325 1125 3355
rect 1155 3325 1160 3355
rect 840 3320 1160 3325
rect -80 3275 0 3280
rect -80 3245 -75 3275
rect -45 3245 0 3275
rect -80 3240 0 3245
rect -80 3195 0 3200
rect -80 3165 -75 3195
rect -45 3165 0 3195
rect -80 3160 0 3165
rect -240 3115 0 3120
rect -240 3085 -235 3115
rect -205 3085 0 3115
rect -240 3080 0 3085
rect -240 3035 0 3040
rect -240 3005 -235 3035
rect -205 3005 0 3035
rect -240 3000 0 3005
rect -80 2955 0 2960
rect -80 2925 -75 2955
rect -45 2925 0 2955
rect -80 2920 0 2925
rect -80 2875 0 2880
rect -80 2845 -75 2875
rect -45 2845 0 2875
rect -80 2840 0 2845
rect -80 2595 0 2600
rect -80 2565 -75 2595
rect -45 2565 0 2595
rect -80 2560 0 2565
rect 840 2515 920 2520
rect 840 2485 885 2515
rect 915 2485 920 2515
rect 840 2480 920 2485
rect 840 2435 1000 2440
rect 840 2405 965 2435
rect 995 2405 1000 2435
rect 840 2400 1000 2405
rect 840 2355 1080 2360
rect 840 2325 1045 2355
rect 1075 2325 1080 2355
rect 840 2320 1080 2325
rect 840 2275 1160 2280
rect 840 2245 1125 2275
rect 1155 2245 1160 2275
rect 840 2240 1160 2245
rect -80 2195 0 2200
rect -80 2165 -75 2195
rect -45 2165 0 2195
rect -80 2160 0 2165
rect -80 2115 0 2120
rect -80 2085 -75 2115
rect -45 2085 0 2115
rect -80 2080 0 2085
rect -320 2035 0 2040
rect -320 2005 -315 2035
rect -285 2005 0 2035
rect -320 2000 0 2005
rect -400 1955 0 1960
rect -400 1925 -395 1955
rect -365 1925 0 1955
rect -400 1920 0 1925
rect -160 1875 0 1880
rect -160 1845 -155 1875
rect -125 1845 0 1875
rect -160 1840 0 1845
rect -80 1795 0 1800
rect -80 1765 -75 1795
rect -45 1765 0 1795
rect -80 1760 0 1765
rect -80 1515 0 1520
rect -80 1485 -75 1515
rect -45 1485 0 1515
rect -80 1480 0 1485
rect 840 1435 1240 1440
rect 840 1405 1205 1435
rect 1235 1405 1240 1435
rect 840 1400 1240 1405
rect 840 1355 1320 1360
rect 840 1325 1285 1355
rect 1315 1325 1320 1355
rect 840 1320 1320 1325
rect 840 1275 1400 1280
rect 840 1245 1365 1275
rect 1395 1245 1400 1275
rect 840 1240 1400 1245
rect 840 1195 1480 1200
rect 840 1165 1445 1195
rect 1475 1165 1480 1195
rect 840 1160 1480 1165
rect -80 1115 0 1120
rect -80 1085 -75 1115
rect -45 1085 0 1115
rect -80 1080 0 1085
rect -80 1035 0 1040
rect -80 1005 -75 1035
rect -45 1005 0 1035
rect -80 1000 0 1005
rect -160 955 0 960
rect -160 925 -155 955
rect -125 925 0 955
rect -160 920 0 925
rect -240 875 0 880
rect -240 845 -235 875
rect -205 845 0 875
rect -240 840 0 845
rect -80 795 0 800
rect -80 765 -75 795
rect -45 765 0 795
rect -80 760 0 765
rect -80 715 0 720
rect -80 685 -75 715
rect -45 685 0 715
rect -80 680 0 685
rect -80 435 0 440
rect -80 405 -75 435
rect -45 405 0 435
rect -80 400 0 405
rect 840 355 1240 360
rect 840 325 1205 355
rect 1235 325 1240 355
rect 840 320 1240 325
rect 840 275 1320 280
rect 840 245 1285 275
rect 1315 245 1320 275
rect 840 240 1320 245
rect 840 195 1400 200
rect 840 165 1365 195
rect 1395 165 1400 195
rect 840 160 1400 165
rect 840 115 1480 120
rect 840 85 1445 115
rect 1475 85 1480 115
rect 840 80 1480 85
rect -80 35 0 40
rect -80 5 -75 35
rect -45 5 0 35
rect -80 0 0 5
rect -400 -45 -360 -40
rect -400 -75 -395 -45
rect -365 -75 -360 -45
rect -400 -125 -360 -75
rect -400 -155 -395 -125
rect -365 -155 -360 -125
rect -400 -160 -360 -155
rect -320 -45 -280 -40
rect -320 -75 -315 -45
rect -285 -75 -280 -45
rect -320 -125 -280 -75
rect -320 -155 -315 -125
rect -285 -155 -280 -125
rect -320 -160 -280 -155
rect 880 -45 920 -40
rect 880 -75 885 -45
rect 915 -75 920 -45
rect 880 -125 920 -75
rect 880 -155 885 -125
rect 915 -155 920 -125
rect 880 -160 920 -155
rect 960 -45 1000 -40
rect 960 -75 965 -45
rect 995 -75 1000 -45
rect 960 -125 1000 -75
rect 960 -155 965 -125
rect 995 -155 1000 -125
rect 960 -160 1000 -155
rect 1040 -45 1080 -40
rect 1040 -75 1045 -45
rect 1075 -75 1080 -45
rect 1040 -125 1080 -75
rect 1040 -155 1045 -125
rect 1075 -155 1080 -125
rect 1040 -160 1080 -155
rect 1120 -45 1160 -40
rect 1120 -75 1125 -45
rect 1155 -75 1160 -45
rect 1120 -125 1160 -75
rect 1120 -155 1125 -125
rect 1155 -155 1160 -125
rect 1120 -160 1160 -155
rect 1200 -45 1240 -40
rect 1200 -75 1205 -45
rect 1235 -75 1240 -45
rect 1200 -125 1240 -75
rect 1200 -155 1205 -125
rect 1235 -155 1240 -125
rect 1200 -160 1240 -155
rect 1280 -45 1320 -40
rect 1280 -75 1285 -45
rect 1315 -75 1320 -45
rect 1280 -125 1320 -75
rect 1280 -155 1285 -125
rect 1315 -155 1320 -125
rect 1280 -160 1320 -155
rect 1360 -45 1400 -40
rect 1360 -75 1365 -45
rect 1395 -75 1400 -45
rect 1360 -125 1400 -75
rect 1360 -155 1365 -125
rect 1395 -155 1400 -125
rect 1360 -160 1400 -155
rect 1440 -45 1480 -40
rect 1440 -75 1445 -45
rect 1475 -75 1480 -45
rect 1440 -125 1480 -75
rect 1440 -155 1445 -125
rect 1475 -155 1480 -125
rect 1440 -160 1480 -155
<< via2 >>
rect -395 4405 -365 4435
rect -395 4325 -365 4355
rect -315 4405 -285 4435
rect -315 4325 -285 4355
rect 885 4405 915 4435
rect 885 4325 915 4355
rect 965 4405 995 4435
rect 965 4325 995 4355
rect 1045 4405 1075 4435
rect 1045 4325 1075 4355
rect 1125 4405 1155 4435
rect 1125 4325 1155 4355
rect 1205 4405 1235 4435
rect 1205 4325 1235 4355
rect 1285 4405 1315 4435
rect 1285 4325 1315 4355
rect 1365 4405 1395 4435
rect 1365 4325 1395 4355
rect 1445 4405 1475 4435
rect 1445 4325 1475 4355
rect -75 4245 -45 4275
rect -395 4165 -365 4195
rect -395 4085 -365 4115
rect -235 4005 -205 4035
rect -75 3925 -45 3955
rect -75 3645 -45 3675
rect 885 3565 915 3595
rect 965 3485 995 3515
rect 1045 3405 1075 3435
rect 1125 3325 1155 3355
rect -75 3245 -45 3275
rect -75 3165 -45 3195
rect -235 3085 -205 3115
rect -235 3005 -205 3035
rect -75 2925 -45 2955
rect -75 2845 -45 2875
rect -75 2565 -45 2595
rect 885 2485 915 2515
rect 965 2405 995 2435
rect 1045 2325 1075 2355
rect 1125 2245 1155 2275
rect -75 2165 -45 2195
rect -75 2085 -45 2115
rect -315 2005 -285 2035
rect -395 1925 -365 1955
rect -155 1845 -125 1875
rect -75 1765 -45 1795
rect -75 1485 -45 1515
rect 1205 1405 1235 1435
rect 1285 1325 1315 1355
rect 1365 1245 1395 1275
rect 1445 1165 1475 1195
rect -75 1085 -45 1115
rect -75 1005 -45 1035
rect -155 925 -125 955
rect -235 845 -205 875
rect -75 765 -45 795
rect -75 685 -45 715
rect -75 405 -45 435
rect 1205 325 1235 355
rect 1285 245 1315 275
rect 1365 165 1395 195
rect 1445 85 1475 115
rect -75 5 -45 35
rect -395 -75 -365 -45
rect -395 -155 -365 -125
rect -315 -75 -285 -45
rect -315 -155 -285 -125
rect 885 -75 915 -45
rect 885 -155 915 -125
rect 965 -75 995 -45
rect 965 -155 995 -125
rect 1045 -75 1075 -45
rect 1045 -155 1075 -125
rect 1125 -75 1155 -45
rect 1125 -155 1155 -125
rect 1205 -75 1235 -45
rect 1205 -155 1235 -125
rect 1285 -75 1315 -45
rect 1285 -155 1315 -125
rect 1365 -75 1395 -45
rect 1365 -155 1395 -125
rect 1445 -75 1475 -45
rect 1445 -155 1475 -125
<< metal3 >>
rect -400 4435 -360 4480
rect -400 4405 -395 4435
rect -365 4405 -360 4435
rect -400 4400 -360 4405
rect -320 4435 -280 4480
rect -320 4405 -315 4435
rect -285 4405 -280 4435
rect -320 4400 -280 4405
rect -400 4355 -360 4360
rect -400 4325 -395 4355
rect -365 4325 -360 4355
rect -400 4195 -360 4325
rect -400 4165 -395 4195
rect -365 4165 -360 4195
rect -400 4115 -360 4165
rect -400 4085 -395 4115
rect -365 4085 -360 4115
rect -400 1955 -360 4085
rect -400 1925 -395 1955
rect -365 1925 -360 1955
rect -400 -45 -360 1925
rect -400 -75 -395 -45
rect -365 -75 -360 -45
rect -400 -80 -360 -75
rect -320 4355 -280 4360
rect -320 4325 -315 4355
rect -285 4325 -280 4355
rect -320 2035 -280 4325
rect -320 2005 -315 2035
rect -285 2005 -280 2035
rect -320 -45 -280 2005
rect -240 4035 -200 4320
rect -240 4005 -235 4035
rect -205 4005 -200 4035
rect -240 3115 -200 4005
rect -240 3085 -235 3115
rect -205 3085 -200 3115
rect -240 3035 -200 3085
rect -240 3005 -235 3035
rect -205 3005 -200 3035
rect -240 875 -200 3005
rect -240 845 -235 875
rect -205 845 -200 875
rect -240 -40 -200 845
rect -160 1875 -120 4320
rect -160 1845 -155 1875
rect -125 1845 -120 1875
rect -160 955 -120 1845
rect -160 925 -155 955
rect -125 925 -120 955
rect -160 -40 -120 925
rect -80 4275 -40 4480
rect 880 4435 920 4480
rect 880 4405 885 4435
rect 915 4405 920 4435
rect 880 4400 920 4405
rect 960 4435 1000 4480
rect 960 4405 965 4435
rect 995 4405 1000 4435
rect 960 4400 1000 4405
rect 1040 4435 1080 4480
rect 1040 4405 1045 4435
rect 1075 4405 1080 4435
rect 1040 4400 1080 4405
rect 1120 4435 1160 4480
rect 1120 4405 1125 4435
rect 1155 4405 1160 4435
rect 1120 4400 1160 4405
rect 1200 4435 1240 4480
rect 1200 4405 1205 4435
rect 1235 4405 1240 4435
rect 1200 4400 1240 4405
rect 1280 4435 1320 4480
rect 1280 4405 1285 4435
rect 1315 4405 1320 4435
rect 1280 4400 1320 4405
rect 1360 4435 1400 4480
rect 1360 4405 1365 4435
rect 1395 4405 1400 4435
rect 1360 4400 1400 4405
rect 1440 4435 1480 4480
rect 1440 4405 1445 4435
rect 1475 4405 1480 4435
rect 1440 4400 1480 4405
rect -80 4245 -75 4275
rect -45 4245 -40 4275
rect -80 3955 -40 4245
rect -80 3925 -75 3955
rect -45 3925 -40 3955
rect -80 3675 -40 3925
rect -80 3645 -75 3675
rect -45 3645 -40 3675
rect -80 3275 -40 3645
rect -80 3245 -75 3275
rect -45 3245 -40 3275
rect -80 3195 -40 3245
rect -80 3165 -75 3195
rect -45 3165 -40 3195
rect -80 2955 -40 3165
rect -80 2925 -75 2955
rect -45 2925 -40 2955
rect -80 2875 -40 2925
rect -80 2845 -75 2875
rect -45 2845 -40 2875
rect -80 2595 -40 2845
rect -80 2565 -75 2595
rect -45 2565 -40 2595
rect -80 2195 -40 2565
rect -80 2165 -75 2195
rect -45 2165 -40 2195
rect -80 2115 -40 2165
rect -80 2085 -75 2115
rect -45 2085 -40 2115
rect -80 1795 -40 2085
rect -80 1765 -75 1795
rect -45 1765 -40 1795
rect -80 1515 -40 1765
rect -80 1485 -75 1515
rect -45 1485 -40 1515
rect -80 1115 -40 1485
rect -80 1085 -75 1115
rect -45 1085 -40 1115
rect -80 1035 -40 1085
rect -80 1005 -75 1035
rect -45 1005 -40 1035
rect -80 795 -40 1005
rect -80 765 -75 795
rect -45 765 -40 795
rect -80 715 -40 765
rect -80 685 -75 715
rect -45 685 -40 715
rect -80 435 -40 685
rect -80 405 -75 435
rect -45 405 -40 435
rect -80 35 -40 405
rect -80 5 -75 35
rect -45 5 -40 35
rect -320 -75 -315 -45
rect -285 -75 -280 -45
rect -320 -80 -280 -75
rect -400 -125 -360 -120
rect -400 -155 -395 -125
rect -365 -155 -360 -125
rect -400 -200 -360 -155
rect -320 -125 -280 -120
rect -320 -155 -315 -125
rect -285 -155 -280 -125
rect -320 -200 -280 -155
rect -80 -200 -40 5
rect 880 4355 920 4360
rect 880 4325 885 4355
rect 915 4325 920 4355
rect 880 3595 920 4325
rect 880 3565 885 3595
rect 915 3565 920 3595
rect 880 2515 920 3565
rect 880 2485 885 2515
rect 915 2485 920 2515
rect 880 -45 920 2485
rect 880 -75 885 -45
rect 915 -75 920 -45
rect 880 -80 920 -75
rect 960 4355 1000 4360
rect 960 4325 965 4355
rect 995 4325 1000 4355
rect 960 3515 1000 4325
rect 960 3485 965 3515
rect 995 3485 1000 3515
rect 960 2435 1000 3485
rect 960 2405 965 2435
rect 995 2405 1000 2435
rect 960 -45 1000 2405
rect 960 -75 965 -45
rect 995 -75 1000 -45
rect 960 -80 1000 -75
rect 1040 4355 1080 4360
rect 1040 4325 1045 4355
rect 1075 4325 1080 4355
rect 1040 3435 1080 4325
rect 1040 3405 1045 3435
rect 1075 3405 1080 3435
rect 1040 2355 1080 3405
rect 1040 2325 1045 2355
rect 1075 2325 1080 2355
rect 1040 -45 1080 2325
rect 1040 -75 1045 -45
rect 1075 -75 1080 -45
rect 1040 -80 1080 -75
rect 1120 4355 1160 4360
rect 1120 4325 1125 4355
rect 1155 4325 1160 4355
rect 1120 3355 1160 4325
rect 1120 3325 1125 3355
rect 1155 3325 1160 3355
rect 1120 2275 1160 3325
rect 1120 2245 1125 2275
rect 1155 2245 1160 2275
rect 1120 -45 1160 2245
rect 1120 -75 1125 -45
rect 1155 -75 1160 -45
rect 1120 -80 1160 -75
rect 1200 4355 1240 4360
rect 1200 4325 1205 4355
rect 1235 4325 1240 4355
rect 1200 1435 1240 4325
rect 1200 1405 1205 1435
rect 1235 1405 1240 1435
rect 1200 355 1240 1405
rect 1200 325 1205 355
rect 1235 325 1240 355
rect 1200 -45 1240 325
rect 1200 -75 1205 -45
rect 1235 -75 1240 -45
rect 1200 -80 1240 -75
rect 1280 4355 1320 4360
rect 1280 4325 1285 4355
rect 1315 4325 1320 4355
rect 1280 1355 1320 4325
rect 1280 1325 1285 1355
rect 1315 1325 1320 1355
rect 1280 275 1320 1325
rect 1280 245 1285 275
rect 1315 245 1320 275
rect 1280 -45 1320 245
rect 1280 -75 1285 -45
rect 1315 -75 1320 -45
rect 1280 -80 1320 -75
rect 1360 4355 1400 4360
rect 1360 4325 1365 4355
rect 1395 4325 1400 4355
rect 1360 1275 1400 4325
rect 1360 1245 1365 1275
rect 1395 1245 1400 1275
rect 1360 195 1400 1245
rect 1360 165 1365 195
rect 1395 165 1400 195
rect 1360 -45 1400 165
rect 1360 -75 1365 -45
rect 1395 -75 1400 -45
rect 1360 -80 1400 -75
rect 1440 4355 1480 4360
rect 1440 4325 1445 4355
rect 1475 4325 1480 4355
rect 1440 1195 1480 4325
rect 1440 1165 1445 1195
rect 1475 1165 1480 1195
rect 1440 115 1480 1165
rect 1440 85 1445 115
rect 1475 85 1480 115
rect 1440 -45 1480 85
rect 1440 -75 1445 -45
rect 1475 -75 1480 -45
rect 1440 -80 1480 -75
rect 880 -125 920 -120
rect 880 -155 885 -125
rect 915 -155 920 -125
rect 880 -200 920 -155
rect 960 -125 1000 -120
rect 960 -155 965 -125
rect 995 -155 1000 -125
rect 960 -200 1000 -155
rect 1040 -125 1080 -120
rect 1040 -155 1045 -125
rect 1075 -155 1080 -125
rect 1040 -200 1080 -155
rect 1120 -125 1160 -120
rect 1120 -155 1125 -125
rect 1155 -155 1160 -125
rect 1120 -200 1160 -155
rect 1200 -125 1240 -120
rect 1200 -155 1205 -125
rect 1235 -155 1240 -125
rect 1200 -200 1240 -155
rect 1280 -125 1320 -120
rect 1280 -155 1285 -125
rect 1315 -155 1320 -125
rect 1280 -200 1320 -155
rect 1360 -125 1400 -120
rect 1360 -155 1365 -125
rect 1395 -155 1400 -125
rect 1360 -200 1400 -155
rect 1440 -125 1480 -120
rect 1440 -155 1445 -125
rect 1475 -155 1480 -125
rect 1440 -200 1480 -155
use prognmos  prognmos_3
timestamp 1642599340
transform 1 0 120 0 1 2680
box -120 -520 720 520
use prognmos  prognmos_2
timestamp 1642599340
transform 1 0 120 0 1 3760
box -120 -520 720 520
use prognmos  prognmos_1
timestamp 1642599340
transform 1 0 120 0 1 1600
box -120 -520 720 520
use prognmos  prognmos_0
timestamp 1642599340
transform 1 0 120 0 1 520
box -120 -520 720 520
<< labels >>
rlabel metal3 -400 4440 -360 4480 0 ii
port 1 nsew
rlabel metal3 -320 4440 -280 4480 0 io
port 2 nsew
rlabel metal3 -80 4440 -40 4480 0 vss
port 5 nsew
rlabel metal3 880 4440 920 4480 0 a1
port 6 nsew
rlabel metal3 960 4440 1000 4480 0 a2
port 7 nsew
rlabel metal3 1040 4440 1080 4480 0 a3
port 8 nsew
rlabel metal3 1120 4440 1160 4480 0 a4
port 9 nsew
rlabel metal3 1200 4440 1240 4480 0 b1
port 10 nsew
rlabel metal3 1280 4440 1320 4480 0 b2
port 11 nsew
rlabel metal3 1360 4440 1400 4480 0 b3
port 12 nsew
rlabel metal3 1440 4440 1480 4480 0 b4
port 13 nsew
rlabel metal3 -400 -200 -360 -160 0 ii
port 1 nsew
rlabel metal3 -320 -200 -280 -160 0 io
port 2 nsew
rlabel metal3 -80 -200 -40 -160 0 vss
port 5 nsew
rlabel metal3 880 -200 920 -160 0 a1
port 6 nsew
rlabel metal3 960 -200 1000 -160 0 a2
port 7 nsew
rlabel metal3 1040 -200 1080 -160 0 a3
port 8 nsew
rlabel metal3 1120 -200 1160 -160 0 a4
port 9 nsew
rlabel metal3 1200 -200 1240 -160 0 b1
port 10 nsew
rlabel metal3 1280 -200 1320 -160 0 b2
port 11 nsew
rlabel metal3 1360 -200 1400 -160 0 b3
port 12 nsew
rlabel metal3 1440 -200 1480 -160 0 b4
port 13 nsew
rlabel metal3 -240 -40 -200 0 0 xl
rlabel metal3 -160 -40 -120 0 0 xr
<< end >>
